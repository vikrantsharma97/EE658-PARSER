1 1 0 1 0
1 2 0 2 0
1 3 0 1 0
2 4 1 2
2 5 1 2
0 6 7 3 2 1 4
2 7 1 6
2 8 1 5
2 9 1 5
2 10 1 6
2 11 1 6
0 12 2 3 2 7 8
2 13 1 12
2 14 1 12
2 15 1 12
0 16 2 2 2 10 13
0 17 5 1 1 14
2 18 1 16
2 19 1 16
0 20 5 2 1 19
2 21 1 20
2 22 1 20
0 23 2 1 2 9 22
3 24 6 0 2 11 18
3 25 3 0 2 17 21
3 26 6 0 3 3 15 23